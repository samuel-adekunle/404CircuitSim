* C:\users\sam\My Documents\LTspiceXVII\Draft1.asc
R1 N003 0 1
V1 N001 0 5
R2 N003 N001 1
R3 N002 N001 {R}
R4 N002 N003 1
R5 N003 N002 1
V2 N003 N004 5
R6 N004 0 1
.step param R 1 1001 1
.op
.backanno
.end
