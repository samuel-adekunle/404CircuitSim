* C:\users\sam\My Documents\LTspiceXVII\Draft2.asc
I1 0 N001 SINE(0 100m 100)
R1 N002 N001 1k
L1 N002 0 100m
R2 N003 N002 100
L2 N003 0 10m
.tran 0 1 0 0.1m
.backanno
.end
