* C:\users\sam\My Documents\LTspiceXVII\Draft2.asc
R1 N004 N001 1k
L1 N004 0 100m
R2 N005 N004 100
L2 N005 0 10m
I1 0 N001 SINE(0 100m 100)
R3 N002 N001 100
C1 N003 N002 10u
R4 N003 N005 50
I2 N002 N004 SINE(0 100m 100)
.tran 0 0.5 0 0.05m
.backanno
.end